package base_pkg;

    

endpackage