`ifndef _DEPENDENCIES_SVH_
`define _DEPENDENCIES_SVH_

`endif